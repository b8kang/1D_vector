##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 08:14:32 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 460.0000 BY 620.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 307.7500 0.6000 307.8500 ;
    END
  END clk
  PIN sum_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0500 0.0000 20.1500 0.6000 ;
    END
  END sum_out[159]
  PIN sum_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.6500 0.0000 22.7500 0.6000 ;
    END
  END sum_out[158]
  PIN sum_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2500 0.0000 25.3500 0.6000 ;
    END
  END sum_out[157]
  PIN sum_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.8500 0.0000 27.9500 0.6000 ;
    END
  END sum_out[156]
  PIN sum_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.4500 0.0000 30.5500 0.6000 ;
    END
  END sum_out[155]
  PIN sum_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0500 0.0000 33.1500 0.6000 ;
    END
  END sum_out[154]
  PIN sum_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.6500 0.0000 35.7500 0.6000 ;
    END
  END sum_out[153]
  PIN sum_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.2500 0.0000 38.3500 0.6000 ;
    END
  END sum_out[152]
  PIN sum_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8500 0.0000 40.9500 0.6000 ;
    END
  END sum_out[151]
  PIN sum_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.4500 0.0000 43.5500 0.6000 ;
    END
  END sum_out[150]
  PIN sum_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.0500 0.0000 46.1500 0.6000 ;
    END
  END sum_out[149]
  PIN sum_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.6500 0.0000 48.7500 0.6000 ;
    END
  END sum_out[148]
  PIN sum_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.2500 0.0000 51.3500 0.6000 ;
    END
  END sum_out[147]
  PIN sum_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.8500 0.0000 53.9500 0.6000 ;
    END
  END sum_out[146]
  PIN sum_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.4500 0.0000 56.5500 0.6000 ;
    END
  END sum_out[145]
  PIN sum_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.0500 0.0000 59.1500 0.6000 ;
    END
  END sum_out[144]
  PIN sum_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.6500 0.0000 61.7500 0.6000 ;
    END
  END sum_out[143]
  PIN sum_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.2500 0.0000 64.3500 0.6000 ;
    END
  END sum_out[142]
  PIN sum_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 0.0000 66.9500 0.6000 ;
    END
  END sum_out[141]
  PIN sum_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.4500 0.0000 69.5500 0.6000 ;
    END
  END sum_out[140]
  PIN sum_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.0500 0.0000 72.1500 0.6000 ;
    END
  END sum_out[139]
  PIN sum_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.6500 0.0000 74.7500 0.6000 ;
    END
  END sum_out[138]
  PIN sum_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.2500 0.0000 77.3500 0.6000 ;
    END
  END sum_out[137]
  PIN sum_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.8500 0.0000 79.9500 0.6000 ;
    END
  END sum_out[136]
  PIN sum_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.4500 0.0000 82.5500 0.6000 ;
    END
  END sum_out[135]
  PIN sum_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.0500 0.0000 85.1500 0.6000 ;
    END
  END sum_out[134]
  PIN sum_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.6500 0.0000 87.7500 0.6000 ;
    END
  END sum_out[133]
  PIN sum_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.2500 0.0000 90.3500 0.6000 ;
    END
  END sum_out[132]
  PIN sum_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.8500 0.0000 92.9500 0.6000 ;
    END
  END sum_out[131]
  PIN sum_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.4500 0.0000 95.5500 0.6000 ;
    END
  END sum_out[130]
  PIN sum_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 0.0000 98.1500 0.6000 ;
    END
  END sum_out[129]
  PIN sum_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.6500 0.0000 100.7500 0.6000 ;
    END
  END sum_out[128]
  PIN sum_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.2500 0.0000 103.3500 0.6000 ;
    END
  END sum_out[127]
  PIN sum_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.8500 0.0000 105.9500 0.6000 ;
    END
  END sum_out[126]
  PIN sum_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 0.0000 108.5500 0.6000 ;
    END
  END sum_out[125]
  PIN sum_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.0500 0.0000 111.1500 0.6000 ;
    END
  END sum_out[124]
  PIN sum_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.6500 0.0000 113.7500 0.6000 ;
    END
  END sum_out[123]
  PIN sum_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.2500 0.0000 116.3500 0.6000 ;
    END
  END sum_out[122]
  PIN sum_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 0.0000 118.9500 0.6000 ;
    END
  END sum_out[121]
  PIN sum_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.4500 0.0000 121.5500 0.6000 ;
    END
  END sum_out[120]
  PIN sum_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.0500 0.0000 124.1500 0.6000 ;
    END
  END sum_out[119]
  PIN sum_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.6500 0.0000 126.7500 0.6000 ;
    END
  END sum_out[118]
  PIN sum_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.2500 0.0000 129.3500 0.6000 ;
    END
  END sum_out[117]
  PIN sum_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.8500 0.0000 131.9500 0.6000 ;
    END
  END sum_out[116]
  PIN sum_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.4500 0.0000 134.5500 0.6000 ;
    END
  END sum_out[115]
  PIN sum_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 0.0000 137.1500 0.6000 ;
    END
  END sum_out[114]
  PIN sum_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.6500 0.0000 139.7500 0.6000 ;
    END
  END sum_out[113]
  PIN sum_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.2500 0.0000 142.3500 0.6000 ;
    END
  END sum_out[112]
  PIN sum_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 0.0000 144.9500 0.6000 ;
    END
  END sum_out[111]
  PIN sum_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.4500 0.0000 147.5500 0.6000 ;
    END
  END sum_out[110]
  PIN sum_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.0500 0.0000 150.1500 0.6000 ;
    END
  END sum_out[109]
  PIN sum_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.6500 0.0000 152.7500 0.6000 ;
    END
  END sum_out[108]
  PIN sum_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.2500 0.0000 155.3500 0.6000 ;
    END
  END sum_out[107]
  PIN sum_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.8500 0.0000 157.9500 0.6000 ;
    END
  END sum_out[106]
  PIN sum_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.4500 0.0000 160.5500 0.6000 ;
    END
  END sum_out[105]
  PIN sum_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.0500 0.0000 163.1500 0.6000 ;
    END
  END sum_out[104]
  PIN sum_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.6500 0.0000 165.7500 0.6000 ;
    END
  END sum_out[103]
  PIN sum_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.2500 0.0000 168.3500 0.6000 ;
    END
  END sum_out[102]
  PIN sum_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.8500 0.0000 170.9500 0.6000 ;
    END
  END sum_out[101]
  PIN sum_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.4500 0.0000 173.5500 0.6000 ;
    END
  END sum_out[100]
  PIN sum_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.0500 0.0000 176.1500 0.6000 ;
    END
  END sum_out[99]
  PIN sum_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.6500 0.0000 178.7500 0.6000 ;
    END
  END sum_out[98]
  PIN sum_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.2500 0.0000 181.3500 0.6000 ;
    END
  END sum_out[97]
  PIN sum_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.8500 0.0000 183.9500 0.6000 ;
    END
  END sum_out[96]
  PIN sum_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.4500 0.0000 186.5500 0.6000 ;
    END
  END sum_out[95]
  PIN sum_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.0500 0.0000 189.1500 0.6000 ;
    END
  END sum_out[94]
  PIN sum_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.6500 0.0000 191.7500 0.6000 ;
    END
  END sum_out[93]
  PIN sum_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.2500 0.0000 194.3500 0.6000 ;
    END
  END sum_out[92]
  PIN sum_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.8500 0.0000 196.9500 0.6000 ;
    END
  END sum_out[91]
  PIN sum_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.4500 0.0000 199.5500 0.6000 ;
    END
  END sum_out[90]
  PIN sum_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.0500 0.0000 202.1500 0.6000 ;
    END
  END sum_out[89]
  PIN sum_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.6500 0.0000 204.7500 0.6000 ;
    END
  END sum_out[88]
  PIN sum_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.2500 0.0000 207.3500 0.6000 ;
    END
  END sum_out[87]
  PIN sum_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.8500 0.0000 209.9500 0.6000 ;
    END
  END sum_out[86]
  PIN sum_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.4500 0.0000 212.5500 0.6000 ;
    END
  END sum_out[85]
  PIN sum_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.0500 0.0000 215.1500 0.6000 ;
    END
  END sum_out[84]
  PIN sum_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.6500 0.0000 217.7500 0.6000 ;
    END
  END sum_out[83]
  PIN sum_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.2500 0.0000 220.3500 0.6000 ;
    END
  END sum_out[82]
  PIN sum_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.8500 0.0000 222.9500 0.6000 ;
    END
  END sum_out[81]
  PIN sum_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.4500 0.0000 225.5500 0.6000 ;
    END
  END sum_out[80]
  PIN sum_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.0500 0.0000 228.1500 0.6000 ;
    END
  END sum_out[79]
  PIN sum_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.6500 0.0000 230.7500 0.6000 ;
    END
  END sum_out[78]
  PIN sum_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.2500 0.0000 233.3500 0.6000 ;
    END
  END sum_out[77]
  PIN sum_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.8500 0.0000 235.9500 0.6000 ;
    END
  END sum_out[76]
  PIN sum_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.4500 0.0000 238.5500 0.6000 ;
    END
  END sum_out[75]
  PIN sum_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.0500 0.0000 241.1500 0.6000 ;
    END
  END sum_out[74]
  PIN sum_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.6500 0.0000 243.7500 0.6000 ;
    END
  END sum_out[73]
  PIN sum_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.2500 0.0000 246.3500 0.6000 ;
    END
  END sum_out[72]
  PIN sum_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.8500 0.0000 248.9500 0.6000 ;
    END
  END sum_out[71]
  PIN sum_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.4500 0.0000 251.5500 0.6000 ;
    END
  END sum_out[70]
  PIN sum_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.0500 0.0000 254.1500 0.6000 ;
    END
  END sum_out[69]
  PIN sum_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.6500 0.0000 256.7500 0.6000 ;
    END
  END sum_out[68]
  PIN sum_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.2500 0.0000 259.3500 0.6000 ;
    END
  END sum_out[67]
  PIN sum_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.8500 0.0000 261.9500 0.6000 ;
    END
  END sum_out[66]
  PIN sum_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.4500 0.0000 264.5500 0.6000 ;
    END
  END sum_out[65]
  PIN sum_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.0500 0.0000 267.1500 0.6000 ;
    END
  END sum_out[64]
  PIN sum_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.6500 0.0000 269.7500 0.6000 ;
    END
  END sum_out[63]
  PIN sum_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.2500 0.0000 272.3500 0.6000 ;
    END
  END sum_out[62]
  PIN sum_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.8500 0.0000 274.9500 0.6000 ;
    END
  END sum_out[61]
  PIN sum_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.4500 0.0000 277.5500 0.6000 ;
    END
  END sum_out[60]
  PIN sum_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.0500 0.0000 280.1500 0.6000 ;
    END
  END sum_out[59]
  PIN sum_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.6500 0.0000 282.7500 0.6000 ;
    END
  END sum_out[58]
  PIN sum_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.2500 0.0000 285.3500 0.6000 ;
    END
  END sum_out[57]
  PIN sum_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.8500 0.0000 287.9500 0.6000 ;
    END
  END sum_out[56]
  PIN sum_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.4500 0.0000 290.5500 0.6000 ;
    END
  END sum_out[55]
  PIN sum_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.0500 0.0000 293.1500 0.6000 ;
    END
  END sum_out[54]
  PIN sum_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.6500 0.0000 295.7500 0.6000 ;
    END
  END sum_out[53]
  PIN sum_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.2500 0.0000 298.3500 0.6000 ;
    END
  END sum_out[52]
  PIN sum_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.8500 0.0000 300.9500 0.6000 ;
    END
  END sum_out[51]
  PIN sum_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.4500 0.0000 303.5500 0.6000 ;
    END
  END sum_out[50]
  PIN sum_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.0500 0.0000 306.1500 0.6000 ;
    END
  END sum_out[49]
  PIN sum_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.6500 0.0000 308.7500 0.6000 ;
    END
  END sum_out[48]
  PIN sum_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.2500 0.0000 311.3500 0.6000 ;
    END
  END sum_out[47]
  PIN sum_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.8500 0.0000 313.9500 0.6000 ;
    END
  END sum_out[46]
  PIN sum_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.4500 0.0000 316.5500 0.6000 ;
    END
  END sum_out[45]
  PIN sum_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.0500 0.0000 319.1500 0.6000 ;
    END
  END sum_out[44]
  PIN sum_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.6500 0.0000 321.7500 0.6000 ;
    END
  END sum_out[43]
  PIN sum_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.2500 0.0000 324.3500 0.6000 ;
    END
  END sum_out[42]
  PIN sum_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.8500 0.0000 326.9500 0.6000 ;
    END
  END sum_out[41]
  PIN sum_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.4500 0.0000 329.5500 0.6000 ;
    END
  END sum_out[40]
  PIN sum_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.0500 0.0000 332.1500 0.6000 ;
    END
  END sum_out[39]
  PIN sum_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.6500 0.0000 334.7500 0.6000 ;
    END
  END sum_out[38]
  PIN sum_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.2500 0.0000 337.3500 0.6000 ;
    END
  END sum_out[37]
  PIN sum_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.8500 0.0000 339.9500 0.6000 ;
    END
  END sum_out[36]
  PIN sum_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.4500 0.0000 342.5500 0.6000 ;
    END
  END sum_out[35]
  PIN sum_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.0500 0.0000 345.1500 0.6000 ;
    END
  END sum_out[34]
  PIN sum_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.6500 0.0000 347.7500 0.6000 ;
    END
  END sum_out[33]
  PIN sum_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.2500 0.0000 350.3500 0.6000 ;
    END
  END sum_out[32]
  PIN sum_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.8500 0.0000 352.9500 0.6000 ;
    END
  END sum_out[31]
  PIN sum_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.4500 0.0000 355.5500 0.6000 ;
    END
  END sum_out[30]
  PIN sum_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.0500 0.0000 358.1500 0.6000 ;
    END
  END sum_out[29]
  PIN sum_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.6500 0.0000 360.7500 0.6000 ;
    END
  END sum_out[28]
  PIN sum_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.2500 0.0000 363.3500 0.6000 ;
    END
  END sum_out[27]
  PIN sum_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.8500 0.0000 365.9500 0.6000 ;
    END
  END sum_out[26]
  PIN sum_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.4500 0.0000 368.5500 0.6000 ;
    END
  END sum_out[25]
  PIN sum_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.0500 0.0000 371.1500 0.6000 ;
    END
  END sum_out[24]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.6500 0.0000 373.7500 0.6000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.2500 0.0000 376.3500 0.6000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.8500 0.0000 378.9500 0.6000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.4500 0.0000 381.5500 0.6000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.0500 0.0000 384.1500 0.6000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.6500 0.0000 386.7500 0.6000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.2500 0.0000 389.3500 0.6000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.8500 0.0000 391.9500 0.6000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.4500 0.0000 394.5500 0.6000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.0500 0.0000 397.1500 0.6000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.6500 0.0000 399.7500 0.6000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.2500 0.0000 402.3500 0.6000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.8500 0.0000 404.9500 0.6000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.4500 0.0000 407.5500 0.6000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.0500 0.0000 410.1500 0.6000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.6500 0.0000 412.7500 0.6000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.2500 0.0000 415.3500 0.6000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.8500 0.0000 417.9500 0.6000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.4500 0.0000 420.5500 0.6000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.0500 0.0000 423.1500 0.6000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.6500 0.0000 425.7500 0.6000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.2500 0.0000 428.3500 0.6000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.8500 0.0000 430.9500 0.6000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.4500 0.0000 433.5500 0.6000 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.0500 619.4000 138.1500 620.0000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.0500 619.4000 142.1500 620.0000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.0500 619.4000 146.1500 620.0000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.0500 619.4000 150.1500 620.0000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.0500 619.4000 154.1500 620.0000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.0500 619.4000 158.1500 620.0000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.0500 619.4000 162.1500 620.0000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.0500 619.4000 166.1500 620.0000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.0500 619.4000 170.1500 620.0000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.0500 619.4000 174.1500 620.0000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.0500 619.4000 178.1500 620.0000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.0500 619.4000 182.1500 620.0000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.0500 619.4000 186.1500 620.0000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.0500 619.4000 190.1500 620.0000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.0500 619.4000 194.1500 620.0000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.0500 619.4000 198.1500 620.0000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.0500 619.4000 202.1500 620.0000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.0500 619.4000 206.1500 620.0000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.0500 619.4000 210.1500 620.0000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.0500 619.4000 214.1500 620.0000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.0500 619.4000 218.1500 620.0000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.0500 619.4000 222.1500 620.0000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.0500 619.4000 226.1500 620.0000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.0500 619.4000 230.1500 620.0000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.0500 619.4000 234.1500 620.0000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.0500 619.4000 238.1500 620.0000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.0500 619.4000 242.1500 620.0000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.0500 619.4000 246.1500 620.0000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.0500 619.4000 250.1500 620.0000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.0500 619.4000 254.1500 620.0000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.0500 619.4000 258.1500 620.0000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.0500 619.4000 262.1500 620.0000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.0500 619.4000 266.1500 620.0000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.0500 619.4000 270.1500 620.0000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.0500 619.4000 274.1500 620.0000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.0500 619.4000 278.1500 620.0000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.0500 619.4000 282.1500 620.0000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.0500 619.4000 286.1500 620.0000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.0500 619.4000 290.1500 620.0000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.0500 619.4000 294.1500 620.0000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.0500 619.4000 298.1500 620.0000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.0500 619.4000 302.1500 620.0000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.0500 619.4000 306.1500 620.0000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.0500 619.4000 310.1500 620.0000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.0500 619.4000 314.1500 620.0000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.0500 619.4000 318.1500 620.0000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.0500 619.4000 322.1500 620.0000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.0500 619.4000 326.1500 620.0000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.0500 619.4000 330.1500 620.0000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.0500 619.4000 334.1500 620.0000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.0500 619.4000 338.1500 620.0000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.0500 619.4000 342.1500 620.0000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.0500 619.4000 346.1500 620.0000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.0500 619.4000 350.1500 620.0000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.0500 619.4000 354.1500 620.0000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.0500 619.4000 358.1500 620.0000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.0500 619.4000 362.1500 620.0000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.0500 619.4000 366.1500 620.0000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.0500 619.4000 370.1500 620.0000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.0500 619.4000 374.1500 620.0000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.0500 619.4000 378.1500 620.0000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.0500 619.4000 382.1500 620.0000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.0500 619.4000 386.1500 620.0000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.0500 619.4000 390.1500 620.0000 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 71.1500 460.0000 71.2500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 74.1500 460.0000 74.2500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 77.1500 460.0000 77.2500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 80.1500 460.0000 80.2500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 83.1500 460.0000 83.2500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 86.1500 460.0000 86.2500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 89.1500 460.0000 89.2500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 92.1500 460.0000 92.2500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 95.1500 460.0000 95.2500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 98.1500 460.0000 98.2500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 101.1500 460.0000 101.2500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 104.1500 460.0000 104.2500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 107.1500 460.0000 107.2500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 110.1500 460.0000 110.2500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 113.1500 460.0000 113.2500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 116.1500 460.0000 116.2500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 119.1500 460.0000 119.2500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 122.1500 460.0000 122.2500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 125.1500 460.0000 125.2500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 128.1500 460.0000 128.2500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 131.1500 460.0000 131.2500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 134.1500 460.0000 134.2500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 137.1500 460.0000 137.2500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 140.1500 460.0000 140.2500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 143.1500 460.0000 143.2500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 146.1500 460.0000 146.2500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 149.1500 460.0000 149.2500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 152.1500 460.0000 152.2500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 155.1500 460.0000 155.2500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 158.1500 460.0000 158.2500 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 161.1500 460.0000 161.2500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 164.1500 460.0000 164.2500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 167.1500 460.0000 167.2500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 170.1500 460.0000 170.2500 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 173.1500 460.0000 173.2500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 176.1500 460.0000 176.2500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 179.1500 460.0000 179.2500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 182.1500 460.0000 182.2500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 185.1500 460.0000 185.2500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 188.1500 460.0000 188.2500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 191.1500 460.0000 191.2500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 194.1500 460.0000 194.2500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 197.1500 460.0000 197.2500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 200.1500 460.0000 200.2500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 203.1500 460.0000 203.2500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 206.1500 460.0000 206.2500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 209.1500 460.0000 209.2500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 212.1500 460.0000 212.2500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 215.1500 460.0000 215.2500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 218.1500 460.0000 218.2500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 221.1500 460.0000 221.2500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 224.1500 460.0000 224.2500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 227.1500 460.0000 227.2500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 230.1500 460.0000 230.2500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 233.1500 460.0000 233.2500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 236.1500 460.0000 236.2500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 239.1500 460.0000 239.2500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 242.1500 460.0000 242.2500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 245.1500 460.0000 245.2500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 248.1500 460.0000 248.2500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 251.1500 460.0000 251.2500 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 254.1500 460.0000 254.2500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 257.1500 460.0000 257.2500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 260.1500 460.0000 260.2500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 263.1500 460.0000 263.2500 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 266.1500 460.0000 266.2500 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 269.1500 460.0000 269.2500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 272.1500 460.0000 272.2500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 275.1500 460.0000 275.2500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 278.1500 460.0000 278.2500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 281.1500 460.0000 281.2500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 284.1500 460.0000 284.2500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 287.1500 460.0000 287.2500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 290.1500 460.0000 290.2500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 293.1500 460.0000 293.2500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 296.1500 460.0000 296.2500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 299.1500 460.0000 299.2500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 302.1500 460.0000 302.2500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 305.1500 460.0000 305.2500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 308.1500 460.0000 308.2500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 311.1500 460.0000 311.2500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 314.1500 460.0000 314.2500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 317.1500 460.0000 317.2500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 320.1500 460.0000 320.2500 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 323.1500 460.0000 323.2500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 326.1500 460.0000 326.2500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 329.1500 460.0000 329.2500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 332.1500 460.0000 332.2500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 335.1500 460.0000 335.2500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 338.1500 460.0000 338.2500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 341.1500 460.0000 341.2500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 344.1500 460.0000 344.2500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 347.1500 460.0000 347.2500 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 350.1500 460.0000 350.2500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 353.1500 460.0000 353.2500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 356.1500 460.0000 356.2500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 359.1500 460.0000 359.2500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 362.1500 460.0000 362.2500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 365.1500 460.0000 365.2500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 368.1500 460.0000 368.2500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 371.1500 460.0000 371.2500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 374.1500 460.0000 374.2500 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 377.1500 460.0000 377.2500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 380.1500 460.0000 380.2500 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 383.1500 460.0000 383.2500 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 386.1500 460.0000 386.2500 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 389.1500 460.0000 389.2500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 392.1500 460.0000 392.2500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 395.1500 460.0000 395.2500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 398.1500 460.0000 398.2500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 401.1500 460.0000 401.2500 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 404.1500 460.0000 404.2500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 407.1500 460.0000 407.2500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 410.1500 460.0000 410.2500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 413.1500 460.0000 413.2500 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 416.1500 460.0000 416.2500 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 419.1500 460.0000 419.2500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 422.1500 460.0000 422.2500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 425.1500 460.0000 425.2500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 428.1500 460.0000 428.2500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 431.1500 460.0000 431.2500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 434.1500 460.0000 434.2500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 437.1500 460.0000 437.2500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 440.1500 460.0000 440.2500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 443.1500 460.0000 443.2500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 446.1500 460.0000 446.2500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 449.1500 460.0000 449.2500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 452.1500 460.0000 452.2500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 455.1500 460.0000 455.2500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 458.1500 460.0000 458.2500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 461.1500 460.0000 461.2500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 464.1500 460.0000 464.2500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 467.1500 460.0000 467.2500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 470.1500 460.0000 470.2500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 473.1500 460.0000 473.2500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 476.1500 460.0000 476.2500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 479.1500 460.0000 479.2500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 482.1500 460.0000 482.2500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 485.1500 460.0000 485.2500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 488.1500 460.0000 488.2500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 491.1500 460.0000 491.2500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 494.1500 460.0000 494.2500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 497.1500 460.0000 497.2500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 500.1500 460.0000 500.2500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 503.1500 460.0000 503.2500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 506.1500 460.0000 506.2500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 509.1500 460.0000 509.2500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 512.1500 460.0000 512.2500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 515.1500 460.0000 515.2500 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 518.1500 460.0000 518.2500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 521.1500 460.0000 521.2500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 524.1500 460.0000 524.2500 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 527.1500 460.0000 527.2500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 530.1500 460.0000 530.2500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 533.1500 460.0000 533.2500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 536.1500 460.0000 536.2500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 539.1500 460.0000 539.2500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 542.1500 460.0000 542.2500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 545.1500 460.0000 545.2500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.4000 548.1500 460.0000 548.2500 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.0500 619.4000 70.1500 620.0000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 619.4000 74.1500 620.0000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.0500 619.4000 78.1500 620.0000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.0500 619.4000 82.1500 620.0000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.0500 619.4000 86.1500 620.0000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.0500 619.4000 90.1500 620.0000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 619.4000 94.1500 620.0000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 619.4000 98.1500 620.0000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 619.4000 102.1500 620.0000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 619.4000 106.1500 620.0000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 619.4000 110.1500 620.0000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.0500 619.4000 114.1500 620.0000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.0500 619.4000 118.1500 620.0000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.0500 619.4000 122.1500 620.0000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.0500 619.4000 126.1500 620.0000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.0500 619.4000 130.1500 620.0000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.0500 619.4000 134.1500 620.0000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 311.7500 0.6000 311.8500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 460.0000 620.0000 ;
    LAYER M2 ;
      RECT 390.2500 619.3000 460.0000 620.0000 ;
      RECT 386.2500 619.3000 389.9500 620.0000 ;
      RECT 382.2500 619.3000 385.9500 620.0000 ;
      RECT 378.2500 619.3000 381.9500 620.0000 ;
      RECT 374.2500 619.3000 377.9500 620.0000 ;
      RECT 370.2500 619.3000 373.9500 620.0000 ;
      RECT 366.2500 619.3000 369.9500 620.0000 ;
      RECT 362.2500 619.3000 365.9500 620.0000 ;
      RECT 358.2500 619.3000 361.9500 620.0000 ;
      RECT 354.2500 619.3000 357.9500 620.0000 ;
      RECT 350.2500 619.3000 353.9500 620.0000 ;
      RECT 346.2500 619.3000 349.9500 620.0000 ;
      RECT 342.2500 619.3000 345.9500 620.0000 ;
      RECT 338.2500 619.3000 341.9500 620.0000 ;
      RECT 334.2500 619.3000 337.9500 620.0000 ;
      RECT 330.2500 619.3000 333.9500 620.0000 ;
      RECT 326.2500 619.3000 329.9500 620.0000 ;
      RECT 322.2500 619.3000 325.9500 620.0000 ;
      RECT 318.2500 619.3000 321.9500 620.0000 ;
      RECT 314.2500 619.3000 317.9500 620.0000 ;
      RECT 310.2500 619.3000 313.9500 620.0000 ;
      RECT 306.2500 619.3000 309.9500 620.0000 ;
      RECT 302.2500 619.3000 305.9500 620.0000 ;
      RECT 298.2500 619.3000 301.9500 620.0000 ;
      RECT 294.2500 619.3000 297.9500 620.0000 ;
      RECT 290.2500 619.3000 293.9500 620.0000 ;
      RECT 286.2500 619.3000 289.9500 620.0000 ;
      RECT 282.2500 619.3000 285.9500 620.0000 ;
      RECT 278.2500 619.3000 281.9500 620.0000 ;
      RECT 274.2500 619.3000 277.9500 620.0000 ;
      RECT 270.2500 619.3000 273.9500 620.0000 ;
      RECT 266.2500 619.3000 269.9500 620.0000 ;
      RECT 262.2500 619.3000 265.9500 620.0000 ;
      RECT 258.2500 619.3000 261.9500 620.0000 ;
      RECT 254.2500 619.3000 257.9500 620.0000 ;
      RECT 250.2500 619.3000 253.9500 620.0000 ;
      RECT 246.2500 619.3000 249.9500 620.0000 ;
      RECT 242.2500 619.3000 245.9500 620.0000 ;
      RECT 238.2500 619.3000 241.9500 620.0000 ;
      RECT 234.2500 619.3000 237.9500 620.0000 ;
      RECT 230.2500 619.3000 233.9500 620.0000 ;
      RECT 226.2500 619.3000 229.9500 620.0000 ;
      RECT 222.2500 619.3000 225.9500 620.0000 ;
      RECT 218.2500 619.3000 221.9500 620.0000 ;
      RECT 214.2500 619.3000 217.9500 620.0000 ;
      RECT 210.2500 619.3000 213.9500 620.0000 ;
      RECT 206.2500 619.3000 209.9500 620.0000 ;
      RECT 202.2500 619.3000 205.9500 620.0000 ;
      RECT 198.2500 619.3000 201.9500 620.0000 ;
      RECT 194.2500 619.3000 197.9500 620.0000 ;
      RECT 190.2500 619.3000 193.9500 620.0000 ;
      RECT 186.2500 619.3000 189.9500 620.0000 ;
      RECT 182.2500 619.3000 185.9500 620.0000 ;
      RECT 178.2500 619.3000 181.9500 620.0000 ;
      RECT 174.2500 619.3000 177.9500 620.0000 ;
      RECT 170.2500 619.3000 173.9500 620.0000 ;
      RECT 166.2500 619.3000 169.9500 620.0000 ;
      RECT 162.2500 619.3000 165.9500 620.0000 ;
      RECT 158.2500 619.3000 161.9500 620.0000 ;
      RECT 154.2500 619.3000 157.9500 620.0000 ;
      RECT 150.2500 619.3000 153.9500 620.0000 ;
      RECT 146.2500 619.3000 149.9500 620.0000 ;
      RECT 142.2500 619.3000 145.9500 620.0000 ;
      RECT 138.2500 619.3000 141.9500 620.0000 ;
      RECT 134.2500 619.3000 137.9500 620.0000 ;
      RECT 130.2500 619.3000 133.9500 620.0000 ;
      RECT 126.2500 619.3000 129.9500 620.0000 ;
      RECT 122.2500 619.3000 125.9500 620.0000 ;
      RECT 118.2500 619.3000 121.9500 620.0000 ;
      RECT 114.2500 619.3000 117.9500 620.0000 ;
      RECT 110.2500 619.3000 113.9500 620.0000 ;
      RECT 106.2500 619.3000 109.9500 620.0000 ;
      RECT 102.2500 619.3000 105.9500 620.0000 ;
      RECT 98.2500 619.3000 101.9500 620.0000 ;
      RECT 94.2500 619.3000 97.9500 620.0000 ;
      RECT 90.2500 619.3000 93.9500 620.0000 ;
      RECT 86.2500 619.3000 89.9500 620.0000 ;
      RECT 82.2500 619.3000 85.9500 620.0000 ;
      RECT 78.2500 619.3000 81.9500 620.0000 ;
      RECT 74.2500 619.3000 77.9500 620.0000 ;
      RECT 70.2500 619.3000 73.9500 620.0000 ;
      RECT 0.0000 619.3000 69.9500 620.0000 ;
      RECT 0.0000 0.7000 460.0000 619.3000 ;
      RECT 433.6500 0.0000 460.0000 0.7000 ;
      RECT 431.0500 0.0000 433.3500 0.7000 ;
      RECT 428.4500 0.0000 430.7500 0.7000 ;
      RECT 425.8500 0.0000 428.1500 0.7000 ;
      RECT 423.2500 0.0000 425.5500 0.7000 ;
      RECT 420.6500 0.0000 422.9500 0.7000 ;
      RECT 418.0500 0.0000 420.3500 0.7000 ;
      RECT 415.4500 0.0000 417.7500 0.7000 ;
      RECT 412.8500 0.0000 415.1500 0.7000 ;
      RECT 410.2500 0.0000 412.5500 0.7000 ;
      RECT 407.6500 0.0000 409.9500 0.7000 ;
      RECT 405.0500 0.0000 407.3500 0.7000 ;
      RECT 402.4500 0.0000 404.7500 0.7000 ;
      RECT 399.8500 0.0000 402.1500 0.7000 ;
      RECT 397.2500 0.0000 399.5500 0.7000 ;
      RECT 394.6500 0.0000 396.9500 0.7000 ;
      RECT 392.0500 0.0000 394.3500 0.7000 ;
      RECT 389.4500 0.0000 391.7500 0.7000 ;
      RECT 386.8500 0.0000 389.1500 0.7000 ;
      RECT 384.2500 0.0000 386.5500 0.7000 ;
      RECT 381.6500 0.0000 383.9500 0.7000 ;
      RECT 379.0500 0.0000 381.3500 0.7000 ;
      RECT 376.4500 0.0000 378.7500 0.7000 ;
      RECT 373.8500 0.0000 376.1500 0.7000 ;
      RECT 371.2500 0.0000 373.5500 0.7000 ;
      RECT 368.6500 0.0000 370.9500 0.7000 ;
      RECT 366.0500 0.0000 368.3500 0.7000 ;
      RECT 363.4500 0.0000 365.7500 0.7000 ;
      RECT 360.8500 0.0000 363.1500 0.7000 ;
      RECT 358.2500 0.0000 360.5500 0.7000 ;
      RECT 355.6500 0.0000 357.9500 0.7000 ;
      RECT 353.0500 0.0000 355.3500 0.7000 ;
      RECT 350.4500 0.0000 352.7500 0.7000 ;
      RECT 347.8500 0.0000 350.1500 0.7000 ;
      RECT 345.2500 0.0000 347.5500 0.7000 ;
      RECT 342.6500 0.0000 344.9500 0.7000 ;
      RECT 340.0500 0.0000 342.3500 0.7000 ;
      RECT 337.4500 0.0000 339.7500 0.7000 ;
      RECT 334.8500 0.0000 337.1500 0.7000 ;
      RECT 332.2500 0.0000 334.5500 0.7000 ;
      RECT 329.6500 0.0000 331.9500 0.7000 ;
      RECT 327.0500 0.0000 329.3500 0.7000 ;
      RECT 324.4500 0.0000 326.7500 0.7000 ;
      RECT 321.8500 0.0000 324.1500 0.7000 ;
      RECT 319.2500 0.0000 321.5500 0.7000 ;
      RECT 316.6500 0.0000 318.9500 0.7000 ;
      RECT 314.0500 0.0000 316.3500 0.7000 ;
      RECT 311.4500 0.0000 313.7500 0.7000 ;
      RECT 308.8500 0.0000 311.1500 0.7000 ;
      RECT 306.2500 0.0000 308.5500 0.7000 ;
      RECT 303.6500 0.0000 305.9500 0.7000 ;
      RECT 301.0500 0.0000 303.3500 0.7000 ;
      RECT 298.4500 0.0000 300.7500 0.7000 ;
      RECT 295.8500 0.0000 298.1500 0.7000 ;
      RECT 293.2500 0.0000 295.5500 0.7000 ;
      RECT 290.6500 0.0000 292.9500 0.7000 ;
      RECT 288.0500 0.0000 290.3500 0.7000 ;
      RECT 285.4500 0.0000 287.7500 0.7000 ;
      RECT 282.8500 0.0000 285.1500 0.7000 ;
      RECT 280.2500 0.0000 282.5500 0.7000 ;
      RECT 277.6500 0.0000 279.9500 0.7000 ;
      RECT 275.0500 0.0000 277.3500 0.7000 ;
      RECT 272.4500 0.0000 274.7500 0.7000 ;
      RECT 269.8500 0.0000 272.1500 0.7000 ;
      RECT 267.2500 0.0000 269.5500 0.7000 ;
      RECT 264.6500 0.0000 266.9500 0.7000 ;
      RECT 262.0500 0.0000 264.3500 0.7000 ;
      RECT 259.4500 0.0000 261.7500 0.7000 ;
      RECT 256.8500 0.0000 259.1500 0.7000 ;
      RECT 254.2500 0.0000 256.5500 0.7000 ;
      RECT 251.6500 0.0000 253.9500 0.7000 ;
      RECT 249.0500 0.0000 251.3500 0.7000 ;
      RECT 246.4500 0.0000 248.7500 0.7000 ;
      RECT 243.8500 0.0000 246.1500 0.7000 ;
      RECT 241.2500 0.0000 243.5500 0.7000 ;
      RECT 238.6500 0.0000 240.9500 0.7000 ;
      RECT 236.0500 0.0000 238.3500 0.7000 ;
      RECT 233.4500 0.0000 235.7500 0.7000 ;
      RECT 230.8500 0.0000 233.1500 0.7000 ;
      RECT 228.2500 0.0000 230.5500 0.7000 ;
      RECT 225.6500 0.0000 227.9500 0.7000 ;
      RECT 223.0500 0.0000 225.3500 0.7000 ;
      RECT 220.4500 0.0000 222.7500 0.7000 ;
      RECT 217.8500 0.0000 220.1500 0.7000 ;
      RECT 215.2500 0.0000 217.5500 0.7000 ;
      RECT 212.6500 0.0000 214.9500 0.7000 ;
      RECT 210.0500 0.0000 212.3500 0.7000 ;
      RECT 207.4500 0.0000 209.7500 0.7000 ;
      RECT 204.8500 0.0000 207.1500 0.7000 ;
      RECT 202.2500 0.0000 204.5500 0.7000 ;
      RECT 199.6500 0.0000 201.9500 0.7000 ;
      RECT 197.0500 0.0000 199.3500 0.7000 ;
      RECT 194.4500 0.0000 196.7500 0.7000 ;
      RECT 191.8500 0.0000 194.1500 0.7000 ;
      RECT 189.2500 0.0000 191.5500 0.7000 ;
      RECT 186.6500 0.0000 188.9500 0.7000 ;
      RECT 184.0500 0.0000 186.3500 0.7000 ;
      RECT 181.4500 0.0000 183.7500 0.7000 ;
      RECT 178.8500 0.0000 181.1500 0.7000 ;
      RECT 176.2500 0.0000 178.5500 0.7000 ;
      RECT 173.6500 0.0000 175.9500 0.7000 ;
      RECT 171.0500 0.0000 173.3500 0.7000 ;
      RECT 168.4500 0.0000 170.7500 0.7000 ;
      RECT 165.8500 0.0000 168.1500 0.7000 ;
      RECT 163.2500 0.0000 165.5500 0.7000 ;
      RECT 160.6500 0.0000 162.9500 0.7000 ;
      RECT 158.0500 0.0000 160.3500 0.7000 ;
      RECT 155.4500 0.0000 157.7500 0.7000 ;
      RECT 152.8500 0.0000 155.1500 0.7000 ;
      RECT 150.2500 0.0000 152.5500 0.7000 ;
      RECT 147.6500 0.0000 149.9500 0.7000 ;
      RECT 145.0500 0.0000 147.3500 0.7000 ;
      RECT 142.4500 0.0000 144.7500 0.7000 ;
      RECT 139.8500 0.0000 142.1500 0.7000 ;
      RECT 137.2500 0.0000 139.5500 0.7000 ;
      RECT 134.6500 0.0000 136.9500 0.7000 ;
      RECT 132.0500 0.0000 134.3500 0.7000 ;
      RECT 129.4500 0.0000 131.7500 0.7000 ;
      RECT 126.8500 0.0000 129.1500 0.7000 ;
      RECT 124.2500 0.0000 126.5500 0.7000 ;
      RECT 121.6500 0.0000 123.9500 0.7000 ;
      RECT 119.0500 0.0000 121.3500 0.7000 ;
      RECT 116.4500 0.0000 118.7500 0.7000 ;
      RECT 113.8500 0.0000 116.1500 0.7000 ;
      RECT 111.2500 0.0000 113.5500 0.7000 ;
      RECT 108.6500 0.0000 110.9500 0.7000 ;
      RECT 106.0500 0.0000 108.3500 0.7000 ;
      RECT 103.4500 0.0000 105.7500 0.7000 ;
      RECT 100.8500 0.0000 103.1500 0.7000 ;
      RECT 98.2500 0.0000 100.5500 0.7000 ;
      RECT 95.6500 0.0000 97.9500 0.7000 ;
      RECT 93.0500 0.0000 95.3500 0.7000 ;
      RECT 90.4500 0.0000 92.7500 0.7000 ;
      RECT 87.8500 0.0000 90.1500 0.7000 ;
      RECT 85.2500 0.0000 87.5500 0.7000 ;
      RECT 82.6500 0.0000 84.9500 0.7000 ;
      RECT 80.0500 0.0000 82.3500 0.7000 ;
      RECT 77.4500 0.0000 79.7500 0.7000 ;
      RECT 74.8500 0.0000 77.1500 0.7000 ;
      RECT 72.2500 0.0000 74.5500 0.7000 ;
      RECT 69.6500 0.0000 71.9500 0.7000 ;
      RECT 67.0500 0.0000 69.3500 0.7000 ;
      RECT 64.4500 0.0000 66.7500 0.7000 ;
      RECT 61.8500 0.0000 64.1500 0.7000 ;
      RECT 59.2500 0.0000 61.5500 0.7000 ;
      RECT 56.6500 0.0000 58.9500 0.7000 ;
      RECT 54.0500 0.0000 56.3500 0.7000 ;
      RECT 51.4500 0.0000 53.7500 0.7000 ;
      RECT 48.8500 0.0000 51.1500 0.7000 ;
      RECT 46.2500 0.0000 48.5500 0.7000 ;
      RECT 43.6500 0.0000 45.9500 0.7000 ;
      RECT 41.0500 0.0000 43.3500 0.7000 ;
      RECT 38.4500 0.0000 40.7500 0.7000 ;
      RECT 35.8500 0.0000 38.1500 0.7000 ;
      RECT 33.2500 0.0000 35.5500 0.7000 ;
      RECT 30.6500 0.0000 32.9500 0.7000 ;
      RECT 28.0500 0.0000 30.3500 0.7000 ;
      RECT 25.4500 0.0000 27.7500 0.7000 ;
      RECT 22.8500 0.0000 25.1500 0.7000 ;
      RECT 20.2500 0.0000 22.5500 0.7000 ;
      RECT 0.0000 0.0000 19.9500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 548.3500 460.0000 620.0000 ;
      RECT 0.0000 548.0500 459.3000 548.3500 ;
      RECT 0.0000 545.3500 460.0000 548.0500 ;
      RECT 0.0000 545.0500 459.3000 545.3500 ;
      RECT 0.0000 542.3500 460.0000 545.0500 ;
      RECT 0.0000 542.0500 459.3000 542.3500 ;
      RECT 0.0000 539.3500 460.0000 542.0500 ;
      RECT 0.0000 539.0500 459.3000 539.3500 ;
      RECT 0.0000 536.3500 460.0000 539.0500 ;
      RECT 0.0000 536.0500 459.3000 536.3500 ;
      RECT 0.0000 533.3500 460.0000 536.0500 ;
      RECT 0.0000 533.0500 459.3000 533.3500 ;
      RECT 0.0000 530.3500 460.0000 533.0500 ;
      RECT 0.0000 530.0500 459.3000 530.3500 ;
      RECT 0.0000 527.3500 460.0000 530.0500 ;
      RECT 0.0000 527.0500 459.3000 527.3500 ;
      RECT 0.0000 524.3500 460.0000 527.0500 ;
      RECT 0.0000 524.0500 459.3000 524.3500 ;
      RECT 0.0000 521.3500 460.0000 524.0500 ;
      RECT 0.0000 521.0500 459.3000 521.3500 ;
      RECT 0.0000 518.3500 460.0000 521.0500 ;
      RECT 0.0000 518.0500 459.3000 518.3500 ;
      RECT 0.0000 515.3500 460.0000 518.0500 ;
      RECT 0.0000 515.0500 459.3000 515.3500 ;
      RECT 0.0000 512.3500 460.0000 515.0500 ;
      RECT 0.0000 512.0500 459.3000 512.3500 ;
      RECT 0.0000 509.3500 460.0000 512.0500 ;
      RECT 0.0000 509.0500 459.3000 509.3500 ;
      RECT 0.0000 506.3500 460.0000 509.0500 ;
      RECT 0.0000 506.0500 459.3000 506.3500 ;
      RECT 0.0000 503.3500 460.0000 506.0500 ;
      RECT 0.0000 503.0500 459.3000 503.3500 ;
      RECT 0.0000 500.3500 460.0000 503.0500 ;
      RECT 0.0000 500.0500 459.3000 500.3500 ;
      RECT 0.0000 497.3500 460.0000 500.0500 ;
      RECT 0.0000 497.0500 459.3000 497.3500 ;
      RECT 0.0000 494.3500 460.0000 497.0500 ;
      RECT 0.0000 494.0500 459.3000 494.3500 ;
      RECT 0.0000 491.3500 460.0000 494.0500 ;
      RECT 0.0000 491.0500 459.3000 491.3500 ;
      RECT 0.0000 488.3500 460.0000 491.0500 ;
      RECT 0.0000 488.0500 459.3000 488.3500 ;
      RECT 0.0000 485.3500 460.0000 488.0500 ;
      RECT 0.0000 485.0500 459.3000 485.3500 ;
      RECT 0.0000 482.3500 460.0000 485.0500 ;
      RECT 0.0000 482.0500 459.3000 482.3500 ;
      RECT 0.0000 479.3500 460.0000 482.0500 ;
      RECT 0.0000 479.0500 459.3000 479.3500 ;
      RECT 0.0000 476.3500 460.0000 479.0500 ;
      RECT 0.0000 476.0500 459.3000 476.3500 ;
      RECT 0.0000 473.3500 460.0000 476.0500 ;
      RECT 0.0000 473.0500 459.3000 473.3500 ;
      RECT 0.0000 470.3500 460.0000 473.0500 ;
      RECT 0.0000 470.0500 459.3000 470.3500 ;
      RECT 0.0000 467.3500 460.0000 470.0500 ;
      RECT 0.0000 467.0500 459.3000 467.3500 ;
      RECT 0.0000 464.3500 460.0000 467.0500 ;
      RECT 0.0000 464.0500 459.3000 464.3500 ;
      RECT 0.0000 461.3500 460.0000 464.0500 ;
      RECT 0.0000 461.0500 459.3000 461.3500 ;
      RECT 0.0000 458.3500 460.0000 461.0500 ;
      RECT 0.0000 458.0500 459.3000 458.3500 ;
      RECT 0.0000 455.3500 460.0000 458.0500 ;
      RECT 0.0000 455.0500 459.3000 455.3500 ;
      RECT 0.0000 452.3500 460.0000 455.0500 ;
      RECT 0.0000 452.0500 459.3000 452.3500 ;
      RECT 0.0000 449.3500 460.0000 452.0500 ;
      RECT 0.0000 449.0500 459.3000 449.3500 ;
      RECT 0.0000 446.3500 460.0000 449.0500 ;
      RECT 0.0000 446.0500 459.3000 446.3500 ;
      RECT 0.0000 443.3500 460.0000 446.0500 ;
      RECT 0.0000 443.0500 459.3000 443.3500 ;
      RECT 0.0000 440.3500 460.0000 443.0500 ;
      RECT 0.0000 440.0500 459.3000 440.3500 ;
      RECT 0.0000 437.3500 460.0000 440.0500 ;
      RECT 0.0000 437.0500 459.3000 437.3500 ;
      RECT 0.0000 434.3500 460.0000 437.0500 ;
      RECT 0.0000 434.0500 459.3000 434.3500 ;
      RECT 0.0000 431.3500 460.0000 434.0500 ;
      RECT 0.0000 431.0500 459.3000 431.3500 ;
      RECT 0.0000 428.3500 460.0000 431.0500 ;
      RECT 0.0000 428.0500 459.3000 428.3500 ;
      RECT 0.0000 425.3500 460.0000 428.0500 ;
      RECT 0.0000 425.0500 459.3000 425.3500 ;
      RECT 0.0000 422.3500 460.0000 425.0500 ;
      RECT 0.0000 422.0500 459.3000 422.3500 ;
      RECT 0.0000 419.3500 460.0000 422.0500 ;
      RECT 0.0000 419.0500 459.3000 419.3500 ;
      RECT 0.0000 416.3500 460.0000 419.0500 ;
      RECT 0.0000 416.0500 459.3000 416.3500 ;
      RECT 0.0000 413.3500 460.0000 416.0500 ;
      RECT 0.0000 413.0500 459.3000 413.3500 ;
      RECT 0.0000 410.3500 460.0000 413.0500 ;
      RECT 0.0000 410.0500 459.3000 410.3500 ;
      RECT 0.0000 407.3500 460.0000 410.0500 ;
      RECT 0.0000 407.0500 459.3000 407.3500 ;
      RECT 0.0000 404.3500 460.0000 407.0500 ;
      RECT 0.0000 404.0500 459.3000 404.3500 ;
      RECT 0.0000 401.3500 460.0000 404.0500 ;
      RECT 0.0000 401.0500 459.3000 401.3500 ;
      RECT 0.0000 398.3500 460.0000 401.0500 ;
      RECT 0.0000 398.0500 459.3000 398.3500 ;
      RECT 0.0000 395.3500 460.0000 398.0500 ;
      RECT 0.0000 395.0500 459.3000 395.3500 ;
      RECT 0.0000 392.3500 460.0000 395.0500 ;
      RECT 0.0000 392.0500 459.3000 392.3500 ;
      RECT 0.0000 389.3500 460.0000 392.0500 ;
      RECT 0.0000 389.0500 459.3000 389.3500 ;
      RECT 0.0000 386.3500 460.0000 389.0500 ;
      RECT 0.0000 386.0500 459.3000 386.3500 ;
      RECT 0.0000 383.3500 460.0000 386.0500 ;
      RECT 0.0000 383.0500 459.3000 383.3500 ;
      RECT 0.0000 380.3500 460.0000 383.0500 ;
      RECT 0.0000 380.0500 459.3000 380.3500 ;
      RECT 0.0000 377.3500 460.0000 380.0500 ;
      RECT 0.0000 377.0500 459.3000 377.3500 ;
      RECT 0.0000 374.3500 460.0000 377.0500 ;
      RECT 0.0000 374.0500 459.3000 374.3500 ;
      RECT 0.0000 371.3500 460.0000 374.0500 ;
      RECT 0.0000 371.0500 459.3000 371.3500 ;
      RECT 0.0000 368.3500 460.0000 371.0500 ;
      RECT 0.0000 368.0500 459.3000 368.3500 ;
      RECT 0.0000 365.3500 460.0000 368.0500 ;
      RECT 0.0000 365.0500 459.3000 365.3500 ;
      RECT 0.0000 362.3500 460.0000 365.0500 ;
      RECT 0.0000 362.0500 459.3000 362.3500 ;
      RECT 0.0000 359.3500 460.0000 362.0500 ;
      RECT 0.0000 359.0500 459.3000 359.3500 ;
      RECT 0.0000 356.3500 460.0000 359.0500 ;
      RECT 0.0000 356.0500 459.3000 356.3500 ;
      RECT 0.0000 353.3500 460.0000 356.0500 ;
      RECT 0.0000 353.0500 459.3000 353.3500 ;
      RECT 0.0000 350.3500 460.0000 353.0500 ;
      RECT 0.0000 350.0500 459.3000 350.3500 ;
      RECT 0.0000 347.3500 460.0000 350.0500 ;
      RECT 0.0000 347.0500 459.3000 347.3500 ;
      RECT 0.0000 344.3500 460.0000 347.0500 ;
      RECT 0.0000 344.0500 459.3000 344.3500 ;
      RECT 0.0000 341.3500 460.0000 344.0500 ;
      RECT 0.0000 341.0500 459.3000 341.3500 ;
      RECT 0.0000 338.3500 460.0000 341.0500 ;
      RECT 0.0000 338.0500 459.3000 338.3500 ;
      RECT 0.0000 335.3500 460.0000 338.0500 ;
      RECT 0.0000 335.0500 459.3000 335.3500 ;
      RECT 0.0000 332.3500 460.0000 335.0500 ;
      RECT 0.0000 332.0500 459.3000 332.3500 ;
      RECT 0.0000 329.3500 460.0000 332.0500 ;
      RECT 0.0000 329.0500 459.3000 329.3500 ;
      RECT 0.0000 326.3500 460.0000 329.0500 ;
      RECT 0.0000 326.0500 459.3000 326.3500 ;
      RECT 0.0000 323.3500 460.0000 326.0500 ;
      RECT 0.0000 323.0500 459.3000 323.3500 ;
      RECT 0.0000 320.3500 460.0000 323.0500 ;
      RECT 0.0000 320.0500 459.3000 320.3500 ;
      RECT 0.0000 317.3500 460.0000 320.0500 ;
      RECT 0.0000 317.0500 459.3000 317.3500 ;
      RECT 0.0000 314.3500 460.0000 317.0500 ;
      RECT 0.0000 314.0500 459.3000 314.3500 ;
      RECT 0.0000 311.9500 460.0000 314.0500 ;
      RECT 0.7000 311.6500 460.0000 311.9500 ;
      RECT 0.0000 311.3500 460.0000 311.6500 ;
      RECT 0.0000 311.0500 459.3000 311.3500 ;
      RECT 0.0000 308.3500 460.0000 311.0500 ;
      RECT 0.0000 308.0500 459.3000 308.3500 ;
      RECT 0.0000 307.9500 460.0000 308.0500 ;
      RECT 0.7000 307.6500 460.0000 307.9500 ;
      RECT 0.0000 305.3500 460.0000 307.6500 ;
      RECT 0.0000 305.0500 459.3000 305.3500 ;
      RECT 0.0000 302.3500 460.0000 305.0500 ;
      RECT 0.0000 302.0500 459.3000 302.3500 ;
      RECT 0.0000 299.3500 460.0000 302.0500 ;
      RECT 0.0000 299.0500 459.3000 299.3500 ;
      RECT 0.0000 296.3500 460.0000 299.0500 ;
      RECT 0.0000 296.0500 459.3000 296.3500 ;
      RECT 0.0000 293.3500 460.0000 296.0500 ;
      RECT 0.0000 293.0500 459.3000 293.3500 ;
      RECT 0.0000 290.3500 460.0000 293.0500 ;
      RECT 0.0000 290.0500 459.3000 290.3500 ;
      RECT 0.0000 287.3500 460.0000 290.0500 ;
      RECT 0.0000 287.0500 459.3000 287.3500 ;
      RECT 0.0000 284.3500 460.0000 287.0500 ;
      RECT 0.0000 284.0500 459.3000 284.3500 ;
      RECT 0.0000 281.3500 460.0000 284.0500 ;
      RECT 0.0000 281.0500 459.3000 281.3500 ;
      RECT 0.0000 278.3500 460.0000 281.0500 ;
      RECT 0.0000 278.0500 459.3000 278.3500 ;
      RECT 0.0000 275.3500 460.0000 278.0500 ;
      RECT 0.0000 275.0500 459.3000 275.3500 ;
      RECT 0.0000 272.3500 460.0000 275.0500 ;
      RECT 0.0000 272.0500 459.3000 272.3500 ;
      RECT 0.0000 269.3500 460.0000 272.0500 ;
      RECT 0.0000 269.0500 459.3000 269.3500 ;
      RECT 0.0000 266.3500 460.0000 269.0500 ;
      RECT 0.0000 266.0500 459.3000 266.3500 ;
      RECT 0.0000 263.3500 460.0000 266.0500 ;
      RECT 0.0000 263.0500 459.3000 263.3500 ;
      RECT 0.0000 260.3500 460.0000 263.0500 ;
      RECT 0.0000 260.0500 459.3000 260.3500 ;
      RECT 0.0000 257.3500 460.0000 260.0500 ;
      RECT 0.0000 257.0500 459.3000 257.3500 ;
      RECT 0.0000 254.3500 460.0000 257.0500 ;
      RECT 0.0000 254.0500 459.3000 254.3500 ;
      RECT 0.0000 251.3500 460.0000 254.0500 ;
      RECT 0.0000 251.0500 459.3000 251.3500 ;
      RECT 0.0000 248.3500 460.0000 251.0500 ;
      RECT 0.0000 248.0500 459.3000 248.3500 ;
      RECT 0.0000 245.3500 460.0000 248.0500 ;
      RECT 0.0000 245.0500 459.3000 245.3500 ;
      RECT 0.0000 242.3500 460.0000 245.0500 ;
      RECT 0.0000 242.0500 459.3000 242.3500 ;
      RECT 0.0000 239.3500 460.0000 242.0500 ;
      RECT 0.0000 239.0500 459.3000 239.3500 ;
      RECT 0.0000 236.3500 460.0000 239.0500 ;
      RECT 0.0000 236.0500 459.3000 236.3500 ;
      RECT 0.0000 233.3500 460.0000 236.0500 ;
      RECT 0.0000 233.0500 459.3000 233.3500 ;
      RECT 0.0000 230.3500 460.0000 233.0500 ;
      RECT 0.0000 230.0500 459.3000 230.3500 ;
      RECT 0.0000 227.3500 460.0000 230.0500 ;
      RECT 0.0000 227.0500 459.3000 227.3500 ;
      RECT 0.0000 224.3500 460.0000 227.0500 ;
      RECT 0.0000 224.0500 459.3000 224.3500 ;
      RECT 0.0000 221.3500 460.0000 224.0500 ;
      RECT 0.0000 221.0500 459.3000 221.3500 ;
      RECT 0.0000 218.3500 460.0000 221.0500 ;
      RECT 0.0000 218.0500 459.3000 218.3500 ;
      RECT 0.0000 215.3500 460.0000 218.0500 ;
      RECT 0.0000 215.0500 459.3000 215.3500 ;
      RECT 0.0000 212.3500 460.0000 215.0500 ;
      RECT 0.0000 212.0500 459.3000 212.3500 ;
      RECT 0.0000 209.3500 460.0000 212.0500 ;
      RECT 0.0000 209.0500 459.3000 209.3500 ;
      RECT 0.0000 206.3500 460.0000 209.0500 ;
      RECT 0.0000 206.0500 459.3000 206.3500 ;
      RECT 0.0000 203.3500 460.0000 206.0500 ;
      RECT 0.0000 203.0500 459.3000 203.3500 ;
      RECT 0.0000 200.3500 460.0000 203.0500 ;
      RECT 0.0000 200.0500 459.3000 200.3500 ;
      RECT 0.0000 197.3500 460.0000 200.0500 ;
      RECT 0.0000 197.0500 459.3000 197.3500 ;
      RECT 0.0000 194.3500 460.0000 197.0500 ;
      RECT 0.0000 194.0500 459.3000 194.3500 ;
      RECT 0.0000 191.3500 460.0000 194.0500 ;
      RECT 0.0000 191.0500 459.3000 191.3500 ;
      RECT 0.0000 188.3500 460.0000 191.0500 ;
      RECT 0.0000 188.0500 459.3000 188.3500 ;
      RECT 0.0000 185.3500 460.0000 188.0500 ;
      RECT 0.0000 185.0500 459.3000 185.3500 ;
      RECT 0.0000 182.3500 460.0000 185.0500 ;
      RECT 0.0000 182.0500 459.3000 182.3500 ;
      RECT 0.0000 179.3500 460.0000 182.0500 ;
      RECT 0.0000 179.0500 459.3000 179.3500 ;
      RECT 0.0000 176.3500 460.0000 179.0500 ;
      RECT 0.0000 176.0500 459.3000 176.3500 ;
      RECT 0.0000 173.3500 460.0000 176.0500 ;
      RECT 0.0000 173.0500 459.3000 173.3500 ;
      RECT 0.0000 170.3500 460.0000 173.0500 ;
      RECT 0.0000 170.0500 459.3000 170.3500 ;
      RECT 0.0000 167.3500 460.0000 170.0500 ;
      RECT 0.0000 167.0500 459.3000 167.3500 ;
      RECT 0.0000 164.3500 460.0000 167.0500 ;
      RECT 0.0000 164.0500 459.3000 164.3500 ;
      RECT 0.0000 161.3500 460.0000 164.0500 ;
      RECT 0.0000 161.0500 459.3000 161.3500 ;
      RECT 0.0000 158.3500 460.0000 161.0500 ;
      RECT 0.0000 158.0500 459.3000 158.3500 ;
      RECT 0.0000 155.3500 460.0000 158.0500 ;
      RECT 0.0000 155.0500 459.3000 155.3500 ;
      RECT 0.0000 152.3500 460.0000 155.0500 ;
      RECT 0.0000 152.0500 459.3000 152.3500 ;
      RECT 0.0000 149.3500 460.0000 152.0500 ;
      RECT 0.0000 149.0500 459.3000 149.3500 ;
      RECT 0.0000 146.3500 460.0000 149.0500 ;
      RECT 0.0000 146.0500 459.3000 146.3500 ;
      RECT 0.0000 143.3500 460.0000 146.0500 ;
      RECT 0.0000 143.0500 459.3000 143.3500 ;
      RECT 0.0000 140.3500 460.0000 143.0500 ;
      RECT 0.0000 140.0500 459.3000 140.3500 ;
      RECT 0.0000 137.3500 460.0000 140.0500 ;
      RECT 0.0000 137.0500 459.3000 137.3500 ;
      RECT 0.0000 134.3500 460.0000 137.0500 ;
      RECT 0.0000 134.0500 459.3000 134.3500 ;
      RECT 0.0000 131.3500 460.0000 134.0500 ;
      RECT 0.0000 131.0500 459.3000 131.3500 ;
      RECT 0.0000 128.3500 460.0000 131.0500 ;
      RECT 0.0000 128.0500 459.3000 128.3500 ;
      RECT 0.0000 125.3500 460.0000 128.0500 ;
      RECT 0.0000 125.0500 459.3000 125.3500 ;
      RECT 0.0000 122.3500 460.0000 125.0500 ;
      RECT 0.0000 122.0500 459.3000 122.3500 ;
      RECT 0.0000 119.3500 460.0000 122.0500 ;
      RECT 0.0000 119.0500 459.3000 119.3500 ;
      RECT 0.0000 116.3500 460.0000 119.0500 ;
      RECT 0.0000 116.0500 459.3000 116.3500 ;
      RECT 0.0000 113.3500 460.0000 116.0500 ;
      RECT 0.0000 113.0500 459.3000 113.3500 ;
      RECT 0.0000 110.3500 460.0000 113.0500 ;
      RECT 0.0000 110.0500 459.3000 110.3500 ;
      RECT 0.0000 107.3500 460.0000 110.0500 ;
      RECT 0.0000 107.0500 459.3000 107.3500 ;
      RECT 0.0000 104.3500 460.0000 107.0500 ;
      RECT 0.0000 104.0500 459.3000 104.3500 ;
      RECT 0.0000 101.3500 460.0000 104.0500 ;
      RECT 0.0000 101.0500 459.3000 101.3500 ;
      RECT 0.0000 98.3500 460.0000 101.0500 ;
      RECT 0.0000 98.0500 459.3000 98.3500 ;
      RECT 0.0000 95.3500 460.0000 98.0500 ;
      RECT 0.0000 95.0500 459.3000 95.3500 ;
      RECT 0.0000 92.3500 460.0000 95.0500 ;
      RECT 0.0000 92.0500 459.3000 92.3500 ;
      RECT 0.0000 89.3500 460.0000 92.0500 ;
      RECT 0.0000 89.0500 459.3000 89.3500 ;
      RECT 0.0000 86.3500 460.0000 89.0500 ;
      RECT 0.0000 86.0500 459.3000 86.3500 ;
      RECT 0.0000 83.3500 460.0000 86.0500 ;
      RECT 0.0000 83.0500 459.3000 83.3500 ;
      RECT 0.0000 80.3500 460.0000 83.0500 ;
      RECT 0.0000 80.0500 459.3000 80.3500 ;
      RECT 0.0000 77.3500 460.0000 80.0500 ;
      RECT 0.0000 77.0500 459.3000 77.3500 ;
      RECT 0.0000 74.3500 460.0000 77.0500 ;
      RECT 0.0000 74.0500 459.3000 74.3500 ;
      RECT 0.0000 71.3500 460.0000 74.0500 ;
      RECT 0.0000 71.0500 459.3000 71.3500 ;
      RECT 0.0000 0.0000 460.0000 71.0500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 460.0000 620.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 460.0000 620.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 460.0000 620.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 460.0000 620.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 460.0000 620.0000 ;
  END
END core

END LIBRARY
